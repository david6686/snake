module left(headx,heady,direction,hex_d);
input headx;
input heady;
input direction;
output hex_d;
endmodule 