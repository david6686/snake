module snake();

endmodule 